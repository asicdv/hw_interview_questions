// ==================================================================== //
// Copyright (c) 2017, Stephen Henry
// All rights reserved.
//
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions
// are met:
//
// * Redistributions of source code must retain the above copyright
//   notice, this list of conditions and the following disclaimer.
//
// * Redistributions in binary form must reproduce the above copyright
//   notice, this list of conditions and the following disclaimer in
//   the documentation and/or other materials provided with the
//   distribution.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS
// "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT
// LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS
// FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
// COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
// INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
// SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
// HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
// STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED
// OF THE POSSIBILITY OF SUCH DAMAGE.
// ==================================================================== //

`include "libv_pkg.vh"

module carry_chain_brent_kung #(parameter int W = 32) (

   //======================================================================== //
   //                                                                         //
   // Generate/Propagate                                                      //
   //                                                                         //
   //======================================================================== //

   //
     input logic [W-1:0]                          p
   , input logic [W-1:0]                          g

   //======================================================================== //
   //                                                                         //
   // Carry-In                                                                //
   //                                                                         //
   //======================================================================== //
     
   //  
   , output logic [W:0]                           c
);

  // ------------------------------------------------------------------------ //
  //
  generate if (W == 128)
    carry_chain_brent_kung_128 u_cc (p, g, c);
  else if (W == 64)
    carry_chain_brent_kung_64 u_cc (p, g, c);
  else if (W == 32)
    carry_chain_brent_kung_32 u_cc (p, g, c);
  else if (W == 16)
    carry_chain_brent_kung_16 u_cc (p, g, c);
//  else
    // A carry chain for this W is not generated by the build scripts.
    // It is necessary to explicitly modify the CMakeLists.txt file to
    // generate it and modify the above generate statements to
    // instantiate it.
//    initial
//      `libtb2_fatal(("Invalid width for Brent Kung carry chain."));
  endgenerate

endmodule // carry_chain_brent_kung
